module simplified_sha256 #(parameter integer NUM_OF_WORDS = 20)(
 input logic  clk, reset_n, start,
 input logic  [15:0] message_addr, output_addr,
 output logic done, mem_clk, mem_we,
 output logic [15:0] mem_addr,
 output logic [31:0] mem_write_data,
 input logic [31:0] mem_read_data);

// parameter integer K[0:63] = '{
parameter integer K[0:63] = '{
   32'h428a2f98,32'h71374491,32'hb5c0fbcf,32'he9b5dba5,32'h3956c25b,32'h59f111f1,32'h923f82a4,32'hab1c5ed5,
   32'hd807aa98,32'h12835b01,32'h243185be,32'h550c7dc3,32'h72be5d74,32'h80deb1fe,32'h9bdc06a7,32'hc19bf174,
   32'he49b69c1,32'hefbe4786,32'h0fc19dc6,32'h240ca1cc,32'h2de92c6f,32'h4a7484aa,32'h5cb0a9dc,32'h76f988da,
   32'h983e5152,32'ha831c66d,32'hb00327c8,32'hbf597fc7,32'hc6e00bf3,32'hd5a79147,32'h06ca6351,32'h14292967,
   32'h27b70a85,32'h2e1b2138,32'h4d2c6dfc,32'h53380d13,32'h650a7354,32'h766a0abb,32'h81c2c92e,32'h92722c85,
   32'ha2bfe8a1,32'ha81a664b,32'hc24b8b70,32'hc76c51a3,32'hd192e819,32'hd6990624,32'hf40e3585,32'h106aa070,
   32'h19a4c116,32'h1e376c08,32'h2748774c,32'h34b0bcb5,32'h391c0cb3,32'h4ed8aa4a,32'h5b9cca4f,32'h682e6ff3,
   32'h748f82ee,32'h78a5636f,32'h84c87814,32'h8cc70208,32'h90befffa,32'ha4506ceb,32'hbef9a3f7,32'hc67178f2
};

localparam [63:0] MessageSize = NUM_OF_WORDS * 32;
localparam int Remainder = MessageSize % 512;
localparam int NumPadZeros = 512 - Remainder - 1 - 64;
localparam int RemainderWords = NUM_OF_WORDS % 16;
localparam logic EvenFit = Remainder == 0;
localparam [7:0] TotalPaddingWidth = 1 + NumPadZeros + 64;

// FSM state variables
enum logic [2:0] {
  IDLE,
  READ,
  BLOCK,
  COMPUTE,
  WRITE
} state;

typedef logic[31:0] logic32;

// NOTE : Below mentioned frame work is for reference purpose.
// Local variables might not be complete and you might have to add more variables
// or modify these variables. Code below is more as a reference.

// Local variables
logic [31:0] w[64];
logic [31:0] message[20];
logic [31:0] wt;
logic [31:0] h0, h1, h2, h3, h4, h5, h6, h7;
logic [31:0] a, b, c, d, e, f, g, h;
logic [ 7:0] i, j, counter;
logic [15:0] offset; // in word address
logic [ 7:0] num_blocks;

logic        cur_we;
logic [15:0] cur_addr;
logic [31:0] cur_write_data;

logic [512:0] memory_block;
logic [ 7:0] tstep;

logic [5:0] t;
logic32 s0;
logic32 s1;




assign num_blocks = determine_num_blocks(NUM_OF_WORDS);
assign tstep = (i - 1);

// Note : Function defined are for reference purpose. Feel free to add more functions or modify below.
// Function to determine number of blocks in memory to fetch
function automatic logic [15:0] determine_num_blocks(input logic [31:0] num_words);
  logic[31:0] size;
begin
    
    size = 32 * num_words;

    if (EvenFit) begin
      determine_num_blocks = size / 512;
    end
    else begin
      determine_num_blocks = (size / 512) + 1;
    end
end
endfunction

function automatic logic[31:0] memory_block_get_block(input logic[7:0] idx);
    logic[31:0] start_addr;
    logic[31:0] end_addr;
begin
    start_addr = (idx+1) * 32;
    end_addr = idx * 32;


end
endfunction


// SHA256 hash round
function automatic logic [255:0] sha256_op(input logic [31:0] a, logic32 b, logic32 c,
  logic32 d, logic32 e, logic32 f, logic32 g, logic32 h, logic32 w,
                                 input logic [7:0] t);
    logic [31:0] S1, S0, ch, maj, t1, t2; // internal signals
begin
    S1 = rightrotate(e, 6) ^ rightrotate(e, 11) ^ rightrotate(e, 25);
    // Student to add remaning code below
    // Refer to SHA256 discussion slides to get logic for this function
    ch = (e & f) ^ ((~e) & g);
    t1 = ch + S1 + h + K[t] + w;
    S0 = rightrotate(a, 2) ^ rightrotate(a, 13) ^ rightrotate(a, 22);
    maj = (a & b) ^ (a & c) ^ (b & c);
    t2 = maj + S0;
    sha256_op = {t1 + t2, a, b, c, d + t1, e, f, g};
end
endfunction

function automatic logic32 word_expand(input logic[5:0] t);
  logic32 s0, s1;
begin
    s0 = rightrotate(w[t-15], 7) ^ rightrotate(w[t-15], 18) ^ (w[t-15] >> 3);
    s1 = rightrotate(w[t-2], 17) ^ rightrotate(w[t-2],  19) ^ (w[t-2]  >> 10);
    word_expand = w[t-16] + s0 + w[t-7] + s1;
end
endfunction


// Generate request to memory
// for reading from memory to get original message
// for writing final computed has value
assign mem_clk = clk;
assign mem_addr = cur_addr + offset;
assign mem_we = cur_we;
assign mem_write_data = cur_write_data;


// rotate `x` right by `r` bits
function automatic logic [31:0] rightrotate(input logic [31:0] x,
                                  input logic [ 7:0] r);
   rightrotate = (x >> r) | (x << (32 - r));
endfunction



// SHA-256 FSM
// Get a BLOCK from the memory, COMPUTE Hash output using SHA256 function
// and write back hash value back to memory
always_ff @(posedge clk, negedge reset_n)
begin
  if (!reset_n) begin
    state <= IDLE;
  end
  else case (state)
    // Initialize hash values h0 to h7 and a to h, other variables and memory we, address offset, etc
    IDLE: begin
        if(start) begin
        // Student to add rest of the code
            h0 <= 'h6a09e667;
            h1 <= 'hbb67ae85;
            h2 <= 'h3c6ef372;
            h3 <= 'ha54ff53a;
            h4 <= 'h510e527f;
            h5 <= 'h9b05688c;
            h6 <= 'h1f83d9ab;
            h7 <= 'h5be0cd19;

            a  <= 'h6a09e667;
            b  <= 'hbb67ae85;
            c  <= 'h3c6ef372;
            d  <= 'ha54ff53a;
            e  <= 'h510e527f;
            f  <= 'h9b05688c;
            g  <= 'h1f83d9ab;
            h  <= 'h5be0cd19;

            // initialize all the counters
            j <= 'b0;
            i <= 'b0;
            offset <= 'b0;
            counter <= 'b0;

            state <= READ;
        end
    end


    READ: begin
        cur_we <= 0;
        cur_addr <= message_addr;

        if (offset <= NUM_OF_WORDS) begin
            // this is to account for delayed appearance of data on mem_read_data
            if (offset > 0) begin
                message[offset-1] <= mem_read_data;
            end
            offset <= offset + 1;
        end
        else begin
            state <= BLOCK;
        end
    end


    // SHA-256 FSM
    // Get a BLOCK from the memory, COMPUTE Hash output using SHA256 function
    // and write back hash value back to memory
    BLOCK: begin
    // Fetch message in 512-bit block size
    // For each of 512-bit block initiate hash value computation
        // in this case deal with padding
        if (!EvenFit && (j + 1) == NUM_OF_WORDS) begin
            for (integer k = 0; k < RemainderWords; k = k + 1) begin
                memory_block[(k*32) +: 32] <= message[(16*j)+k];
            end
            memory_block[TotalPaddingWidth:0] <= {
                1'b1,
                {NumPadZeros{1'b0}},
                MessageSize
            };
        end
        // in this case just fill memory
        else begin
            for (integer k = 0; k < 16; k = k + 32) begin
                memory_block[(k*32) +: 32] <= message[(16*j)+k];
            end
        end
        state <= COMPUTE;
        i <= 0;
    end

    // For each block compute hash function
    // Go back to BLOCK stage after each block hash computation is completed and if
    // there are still number of message blocks available in memory otherwise
    // move to WRITE stage
    COMPUTE: begin
    // 64 processing rounds steps for 512-bit block
        if (i <= 64) begin
            if (i < 16) begin
                w[i] <= memory_block[i*32 +: 32];
            end
            else begin
                w[i] <= word_expand(i);
            end
            i <= i + 1;
            {a, b, c, d, e, f, g, h} <= sha256_op(a, b, c, d, e, f, g, h, w[i], i);
        end
        else begin
            {h0, h1, h2, h3, h4, h5, h6, h7} <= 
                {h0, h1, h2, h3, h4, h5, h6, h7} + {a, b, c, d, e, f, g, h};
            
            if ((j + 1) < num_blocks) begin
                state <= BLOCK;
                j <= j + 1;
            end
            else begin
                state <= WRITE;
            end
        end

    end

    // h0 to h7 each are 32 bit hashes, which makes up total 256 bit value
    // h0 to h7 after compute stage has final computed hash value
    // write back these h0 to h7 to memory starting from output_addr
    WRITE: begin
        cur_addr <= output_addr + counter;
        case(counter)
            0: cur_write_data <= h0;
            1: cur_write_data <= h1;
            2: cur_write_data <= h2;
            3: cur_write_data <= h3;
            4: cur_write_data <= h4;
            5: cur_write_data <= h5;
            6: cur_write_data <= h6;
            7: cur_write_data <= h7;
            default: $display("Error: default in case");
        endcase

        counter <= counter + 1;
    end


    default: begin
        state <= IDLE;
        // $display("We hit default, this should never happen");
    end

   endcase
  end

// Generate done when SHA256 hash computation has finished and moved to IDLE state
assign done = (state == IDLE);

endmodule
