module simplified_sha256 #(parameter integer NUM_OF_WORDS = 20)(
 input logic  clk, reset_n, start,
 input logic  [15:0] message_addr, output_addr,
 output logic done, mem_clk, mem_we,
 output logic [15:0] mem_addr,
 output logic [31:0] mem_write_data,
 input logic [31:0] mem_read_data);

// parameter integer K[0:63] = '{
parameter integer K[0:63] = '{
   32'h428a2f98,32'h71374491,32'hb5c0fbcf,32'he9b5dba5,32'h3956c25b,32'h59f111f1,32'h923f82a4,32'hab1c5ed5,
   32'hd807aa98,32'h12835b01,32'h243185be,32'h550c7dc3,32'h72be5d74,32'h80deb1fe,32'h9bdc06a7,32'hc19bf174,
   32'he49b69c1,32'hefbe4786,32'h0fc19dc6,32'h240ca1cc,32'h2de92c6f,32'h4a7484aa,32'h5cb0a9dc,32'h76f988da,
   32'h983e5152,32'ha831c66d,32'hb00327c8,32'hbf597fc7,32'hc6e00bf3,32'hd5a79147,32'h06ca6351,32'h14292967,
   32'h27b70a85,32'h2e1b2138,32'h4d2c6dfc,32'h53380d13,32'h650a7354,32'h766a0abb,32'h81c2c92e,32'h92722c85,
   32'ha2bfe8a1,32'ha81a664b,32'hc24b8b70,32'hc76c51a3,32'hd192e819,32'hd6990624,32'hf40e3585,32'h106aa070,
   32'h19a4c116,32'h1e376c08,32'h2748774c,32'h34b0bcb5,32'h391c0cb3,32'h4ed8aa4a,32'h5b9cca4f,32'h682e6ff3,
   32'h748f82ee,32'h78a5636f,32'h84c87814,32'h8cc70208,32'h90befffa,32'ha4506ceb,32'hbef9a3f7,32'hc67178f2
};

localparam [63:0] MessageSize = NUM_OF_WORDS * 32;
localparam int Remainder = MessageSize % 512;
localparam int NumPadZeros = 512 - Remainder - 1 - 64;
localparam int RemainderWords = NUM_OF_WORDS % 16;
localparam logic EvenFit = Remainder == 0;
localparam [63:0] TotalPaddingWidth = 512 - Remainder;
localparam [7:0] num_blocks = 2;

// logic [ 7:0] num_blocks;
// assign num_blocks = determine_num_blocks(NUM_OF_WORDS);


// FSM state variables
enum logic [2:0] {
  IDLE,
  READ,
  BLOCK,
  COMPUTE,
  WRITE
} state;

typedef logic[31:0] logic32;

// NOTE : Below mentioned frame work is for reference purpose.
// Local variables might not be complete and you might have to add more variables
// or modify these variables. Code below is more as a reference.

// Local variables
logic [31:0] w[16];
logic [31:0] message[20];
logic [31:0] h0, h1, h2, h3, h4, h5, h6, h7;
logic [31:0] a, b, c, d, e, f, g, h;
logic [ 7:0] i, counter;
logic j;
logic [15:0] offset; // in word address

// logic        cur_we;
// logic [15:0] cur_addr;
logic [31:0] cur_write_data;

logic [511:0] memory_block;

logic32 s0;
logic32 s1;


// function automatic logic [15:0] determine_num_blocks(input logic [31:0] num_words);
//   logic[31:0] size;
// begin
//     
//     size = 32 * num_words;
// 
//     if (EvenFit) begin
//       determine_num_blocks = size / 512;
//     end
//     else begin
//       determine_num_blocks = (size / 512) + 1;
//     end
// end
// endfunction


// SHA256 hash round
function automatic logic [255:0] sha256_op(input logic [31:0] a, logic32 b, logic32 c,
  logic32 d, logic32 e, logic32 f, logic32 g, logic32 h, logic32 w,
                                 input logic [7:0] t);
    logic [31:0] S1, S0, ch, maj, t1, t2; // internal signals
begin
    S1 = rightrotate(e, 6) ^ rightrotate(e, 11) ^ rightrotate(e, 25);
    // Student to add remaning code below
    // Refer to SHA256 discussion slides to get logic for this function
    ch = (e & f) ^ ((~e) & g);
    t1 = ch + S1 + h + K[t] + w;
    S0 = rightrotate(a, 2) ^ rightrotate(a, 13) ^ rightrotate(a, 22);
    maj = (a & b) ^ (a & c) ^ (b & c);
    t2 = maj + S0;
    sha256_op = {t1 + t2, a, b, c, d + t1, e, f, g};
end
endfunction

function automatic logic32 word_expand(input logic[7:0] t);
  logic32 s0, s1;
begin
    if (t < 16) begin
        word_expand = memory_block[t*32 +: 32];
    end
    else begin
        s0 = rightrotate(w[1],7)^rightrotate(w[1],18)^(w[1]>>3);
        s1 = rightrotate(w[14],17)^rightrotate(w[14],19)^(w[14]>>10);
        word_expand = w[0] + s0 + w[9] + s1;
    end
end
endfunction


// Generate request to memory
// for reading from memory to get original message
// for writing final computed has value
assign mem_clk = clk;
// assign mem_addr = cur_addr + offset;
assign mem_addr = (state == WRITE) ? (output_addr + offset) : (message_addr + offset);
assign mem_we = (state == WRITE);
assign mem_write_data = cur_write_data;


// rotate `x` right by `r` bits
function automatic logic [31:0] rightrotate(input logic [31:0] x,
                                  input logic [ 7:0] r);
   rightrotate = (x >> r) | (x << (32 - r));
endfunction


// SHA-256 FSM
// Get a BLOCK from the memory, COMPUTE Hash output using SHA256 function
// and write back hash value back to memory
always_ff @(posedge clk, negedge reset_n)
begin
  if (!reset_n) begin
    state <= IDLE;
  end
  else case (state)
    // Initialize hash values h0 to h7 and a to h, other variables and memory we, address offset, etc
    IDLE: begin
        if(start) begin
$display("TotalPaddingWidth = %d", TotalPaddingWidth);
        // Student to add rest of the code
            h0 <= 'h6a09e667;
            h1 <= 'hbb67ae85;
            h2 <= 'h3c6ef372;
            h3 <= 'ha54ff53a;
            h4 <= 'h510e527f;
            h5 <= 'h9b05688c;
            h6 <= 'h1f83d9ab;
            h7 <= 'h5be0cd19;

            // a  <= 'h6a09e667;
            // b  <= 'hbb67ae85;
            // c  <= 'h3c6ef372;
            // d  <= 'ha54ff53a;
            // e  <= 'h510e527f;
            // f  <= 'h9b05688c;
            // g  <= 'h1f83d9ab;
            // h  <= 'h5be0cd19;

            // initialize all the counters
            j <= 'b0;
            i <= 'b0;
            counter <= 'b0;

            // prep for transition to READ_WAIT
            // state <= READ_WAIT;
            state <= READ;
            offset <= 'b0;
            //cur_we <= 0;
            // cur_addr <= message_addr;

            // $display("NUM_OF_WORDS=%d", NUM_OF_WORDS);
        end
    end


    READ: begin
        if (offset <= NUM_OF_WORDS) begin
            // this is to account for delayed appearance of data on mem_read_data
            if (offset > 0) begin
                message[offset-1] <= mem_read_data;
            end
            offset <= offset + 1;
        end
        else begin
            state <= BLOCK;
        end
    end


    // SHA-256 FSM
    // Get a BLOCK from the memory, COMPUTE Hash output using SHA256 function
    // and write back hash value back to memory
    BLOCK: begin
    // Fetch message in 512-bit block size
    // For each of 512-bit block initiate hash value computation
        // in this case deal with padding
        // if ((j + 1) == num_blocks) begin
        if (j == 1) begin
            // $display("padding");
            for (integer k = 0; k < RemainderWords; k = k + 1) begin
                // memory_block[(k*32) +: 32] <= message[(16*j)+k];
                memory_block[(k*32) +: 32] <= message[16+k];
            end

            // memory_block[511 -: 64] <= MessageSize;
            // memory_block[(511 - 64) -: NumPadZeros] <= {NumPadZeros{1'b0}};
            // memory_block[(511 - 64 - NumPadZeros)] <= 1'b1;
            memory_block[511 -: TotalPaddingWidth] <= {
                // i do not know why we need to multiply size by 2
                // but otherwise it doesn't match the testbench padding
                MessageSize*2,
                {NumPadZeros{1'b0}},
                32'h80000000
            };
        end
        // in this case just fill memory
        else begin
            // $display("not padding");
            for (integer k = 0; k < 16; k = k + 1) begin
                // memory_block[(k*32) +: 32] <= message[(16*j)+k];
                memory_block[(k*32) +: 32] <= message[k];
            end
        end

        // initialize state variables
        a  <= h0;
        b  <= h1;
        c  <= h2;
        d  <= h3;
        e  <= h4;
        f  <= h5;
        g  <= h6;
        h  <= h7;
        state <= COMPUTE;
        i <= 0;
    end

    // For each block compute hash function
    // Go back to BLOCK stage after each block hash computation is completed and if
    // there are still number of message blocks available in memory otherwise
    // move to WRITE stage
    COMPUTE: begin
    // 64 processing rounds steps for 512-bit block
        // if (i == 0) begin
        //     $display("starting COMPUTE");
        //     $display("j = %d, memory_block = %x", j, memory_block);
        //     $display("i = %d", i);
        //     $display("initial a-h state: %p", {a, b, c, d, e, f, g, h});
        // end

        if (i < 64) begin
            w[15] <= word_expand(i);
            for (int n = 0; n < 15; n++) w[n] <= w[n+1];
            i    <= i + 1;
            // $display("real %d: %p", i, sha256_op(a, b, c, d, e, f, g, h, word_expand(i), i));
            {a, b, c, d, e, f, g, h} <= sha256_op(a, b, c, d, e, f, g, h, word_expand(i), i);
        end
        else begin
            // $display("w = %p", w);
            h0 <= h0 + a;
            h1 <= h1 + b;
            h2 <= h2 + c;
            h3 <= h3 + d;
            h4 <= h4 + e;
            h5 <= h5 + f;
            h6 <= h6 + g;
            h7 <= h7 + h;

            if (j == 0) begin
                state <= BLOCK;
                j <= 'b1;
            end
            else begin
                // cur_addr <= output_addr;
                // ugh
                cur_write_data <= h0 + a;
                // cur_we <= 1;
                offset <= 0;
                counter <= 1;
                state  <= WRITE;
            end
        end

    end

    // h0 to h7 each are 32 bit hashes, which makes up total 256 bit value
    // h0 to h7 after compute stage has final computed hash value
    // write back these h0 to h7 to memory starting from output_addr
    WRITE: begin
        case(counter)
            1: cur_write_data <= h1;
            2: cur_write_data <= h2;
            3: cur_write_data <= h3;
            4: cur_write_data <= h4;
            5: cur_write_data <= h5;
            6: cur_write_data <= h6;
            7: cur_write_data <= h7;
            8: state <= IDLE;
            default: $display("Error: default in case");
        endcase

        offset <= offset + 1;
        counter <= counter + 1;
    end


    default: begin
        state <= IDLE;
        // $display("We hit default, this should never happen");
    end

   endcase
  end

// Generate done when SHA256 hash computation has finished and moved to IDLE state
assign done = (state == IDLE);

endmodule
